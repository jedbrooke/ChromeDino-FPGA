//Module for calculating Res = A*B
//Where A,B and C are 4 by 4 matrices.
module Mat_mult(A,B,M);

    //input and output ports.
    //The size 128 bits which is 4*4=16 elements,each of which is 8 bits wide.    
    input wire [127:0] A;
    input wire [127:0] B;
    output wire [127:0] M;
    //internal variables    
    /*reg [127:0] Res;
    reg [7:0] A1 [0:3][0:3];
    reg [7:0] B1 [0:3][0:3];
    reg [7:0] Res1 [0:3][0:3]; 
    integer i,j,k;*/
	 reg [7:0] Res1 [0:3][0:3];
    /*always@ (A or B)
    begin
    //Initialize the matrices-convert 1 D to 3D arrays
        {A1[0][0],A1[0][1],A1[0][2],A1[0][3],A1[1][0],A1[1][1],A1[1][2],A1[1][3],A1[2][0],A1[2][1],A1[2][2],A1[2][3],A1[3][0],A1[3][1],A1[3][2],A1[3][3]} = A;
        {B1[0][0],B1[0][1],B1[0][2],B1[0][3],B1[1][0],B1[1][1],B1[1][2],B1[1][3],B1[2][0],B1[2][1],B1[2][2],B1[2][3],B1[3][0],B1[3][1],B1[3][2],B1[3][3]} = B;
        i = 0;
        j = 0;
        k = 0;
        {Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3]} = 128'd0; //initiBlize to zeros.
        //MRestrix multiplication
        for(i=0;i < 4;i=i+1)
            for(j=0;j < 4;j=j+1)
                for(k=0;k < 4;k=k+1)
                    Res1[i][j] = Res1[i][j] + (A1[i][k] * B1[k][j]);
        //final output assignment - 3D array to 1D array conversion.            
        Res = {Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3]};            
		  
	 end */
	assign M[127:120] = (A[127:120] * B[127:120]) + (A[119:112] * B[95:88]) + (A[111:104] * B[63:56]) + (A[103:96] * B[31:24]);
	assign M[119:112] = (A[127:120] * B[119:112]) + (A[119:112] * B[87:80]) + (A[111:104] * B[55:48]) + (A[103:96] * B[23:16]);
	assign M[111:104] = (A[127:120] * B[111:104]) + (A[119:112] * B[79:72]) + (A[111:104] * B[47:40]) + (A[103:96] * B[15:8]);
	assign M[103:96] = (A[127:120] * B[103:96]) + (A[119:112] * B[71:64]) + (A[111:104] * B[39:32]) + (A[103:96] * B[7:0]);
	assign M[95:88] = (A[95:88] * B[127:120]) + (A[87:80] * B[95:88]) + (A[79:72] * B[63:56]) + (A[71:64] * B[31:24]);
	assign M[87:80] = (A[95:88] * B[119:112]) + (A[87:80] * B[87:80]) + (A[79:72] * B[55:48]) + (A[71:64] * B[23:16]);
	assign M[79:72] = (A[95:88] * B[111:104]) + (A[87:80] * B[79:72]) + (A[79:72] * B[47:40]) + (A[71:64] * B[15:8]);
	assign M[71:64] = (A[95:88] * B[103:96]) + (A[87:80] * B[71:64]) + (A[79:72] * B[39:32]) + (A[71:64] * B[7:0]);
	assign M[63:56] = (A[63:56] * B[127:120]) + (A[55:48] * B[95:88]) + (A[47:40] * B[63:56]) + (A[39:32] * B[31:24]);
	assign M[55:48] = (A[63:56] * B[119:112]) + (A[55:48] * B[87:80]) + (A[47:40] * B[55:48]) + (A[39:32] * B[23:16]);
	assign M[47:40] = (A[63:56] * B[111:104]) + (A[55:48] * B[79:72]) + (A[47:40] * B[47:40]) + (A[39:32] * B[15:8]);
	assign M[39:32] = (A[63:56] * B[103:96]) + (A[55:48] * B[71:64]) + (A[47:40] * B[39:32]) + (A[39:32] * B[7:0]);
	assign M[31:24] = (A[31:24] * B[127:120]) + (A[23:16] * B[95:88]) + (A[15:8] * B[63:56]) + (A[7:0] * B[31:24]);
	assign M[23:16] = (A[31:24] * B[119:112]) + (A[23:16] * B[87:80]) + (A[15:8] * B[55:48]) + (A[7:0] * B[23:16]);
	assign M[15:8] = (A[31:24] * B[111:104]) + (A[23:16] * B[79:72]) + (A[15:8] * B[47:40]) + (A[7:0] * B[15:8]);
	assign M[7:0] = (A[31:24] * B[103:96]) + (A[23:16] * B[71:64]) + (A[15:8] * B[39:32]) + (A[7:0] * B[7:0]);

	always @(*) begin
		{Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3]} = M;
	end

endmodule